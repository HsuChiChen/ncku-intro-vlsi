/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2021 Spring ---------------------- //
// ---------------------- Editor: Tseng Hsin-Yu (Sylvia) --------- //
// ---------------------- Version : v.1.00  ---------------------- //
// ---------------------- Date : 2021.02    ---------------------- //
// ---------------------- priority encoder  ---------------------- // 
/////////////////////////////////////////////////////////////////////

// Module name and I/O port
module encoder(I3,I2,I1,I0,O1,O0);

// Input and output ports declaration
input I3,I2,I1,I0;
output O1,O0;
 
/********* your code ***********/
wire i2,i3,A,B;
not (i2,I2);
not (i3,I3);
and (A,I1,i2,i3);
and (B,I2,i3);
or (O0,A,I3);
or (O1,B,I3);
/******************************/

endmodule
