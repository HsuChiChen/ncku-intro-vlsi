// Don't modify the following code
`define DATA_BITS 9
`define ADDR_BITS 18
`define MEM_SIZE  (1 << `ADDR_BITS)
`define width 256
`define size  256*256

// Add your define below

