/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2021 Spring ---------------------- //
// ---------------------- Editor: Tseng Hsin-Yu (Sylvia) --------- //
// ---------------------- Version : v.1.00  ---------------------- //
// ---------------------- Date : 2021.02    ---------------------- //
// ---------------------- FullAdder  ----------------------------- // 
/////////////////////////////////////////////////////////////////////
// Module name and I/O port
module FullAdder(A,B,Cin,S,Cout);

// Input and output ports declaration
input A,B,Cin;
output S,Cout;

/********* your code ***********/
wire X,Y,Z;
xor (X,A,B);
and (Z,A,B);
and (Y,X,Cin);
xor (S,X,Cin);
or (Cout,Y,Z);
/******************************/

endmodule
