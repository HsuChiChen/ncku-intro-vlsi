/////////////////////////////////////////////////////////////////////
// ---------------------- IVCAD 2021 Spring ---------------------- //
// ---------------------- Editor : Michael  ---------------------- //
// ---------------------- Version : v.1.00  ---------------------- //
// ---------------------- Date : 2021.02.19 ---------------------- //
// ----------------------  Parametric ReLU  ---------------------- //
/////////////////////////////////////////////////////////////////////


module PRelu(in,out);
				
// ---------------------- input  ---------------------- //
input  signed	[`Pixel_DataSize*2:0]	in;
// ---------------------- output ---------------------- //
output  signed	[`Pixel_DataSize*2:0]	out;
// ----------------------  reg   ---------------------- //


// ---------------------- Write down Your design below  ---------------------- //
assign out = (in[`Pixel_DataSize*2] == 1'b1)? $signed(in) >>> 6 : in;


endmodule
